CircuitMaker Text
5.6
Probes: 1
q1[p]
Transient Analysis
0 541 198 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
9961490 0
0
6 Title:
5 Name:
0
0
0
10
11 Resistor:A~
219 144 160 0 2 5
0 6 7
0
0 0 864 90
2 11
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
41290.9 9
0
11 Resistor:A~
219 105 39 0 2 5
0 3 5
0
0 0 864 90
2 3k
-23 3 -9 11
2 R2
-22 -11 -8 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
41290.9 8
0
11 Resistor:A~
219 144 222 0 3 5
0 2 6 -1
0
0 0 864 90
2 1k
9 2 23 10
2 Rl
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
41290.9 7
0
11 Resistor:A~
219 52 69 0 2 5
0 3 4
0
0 0 864 90
2 3k
-24 3 -10 11
2 R3
-22 -11 -8 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
41290.9 6
0
8 Battery~
219 220 105 0 2 5
0 5 2
0
0 0 864 0
3 12V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5283 0 0
2
41290.9 5
0
7 Ground~
168 220 266 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6874 0 0
2
41290.9 4
0
12 NPN Trans:B~
219 139 102 0 3 7
0 5 3 7
0
0 0 832 0
6 BC547A
12 0 54 8
2 Q1
13 -9 27 -1
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
5305 0 0
2
41290.9 3
0
12 SPST Switch~
165 53 224 0 2 11
0 2 3
0
0 0 4704 270
0
2 S1
11 -5 25 3
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
34 0 0
2
41290.9 2
0
12 NPN Trans:B~
219 114 134 0 3 7
0 3 7 6
0
0 0 832 512
6 BC547A
-56 3 -14 11
2 Q2
-55 -8 -41 0
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
969 0 0
2
41290.9 1
0
4 LED~
171 52 33 0 1 2
10 5
0
0 0 864 0
4 LED1
-42 -1 -14 7
2 D1
-41 -12 -27 -4
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8402 0 0
2
41290.9 0
0
15
1 0 3 0 0 16 0 2 0 0 7 2
105 57
105 102
2 2 4 0 0 16 0 10 4 0 0 2
52 43
52 51
1 0 3 0 0 16 0 4 0 0 10 2
52 87
52 102
1 0 5 0 0 16 0 10 0 0 13 3
52 23
52 9
105 9
0 3 6 0 0 16 0 0 9 8 0 3
144 188
105 188
105 152
0 2 7 0 0 16 0 0 9 14 0 3
144 133
144 134
128 134
1 0 3 0 0 16 0 9 0 0 10 2
105 116
105 102
2 1 6 0 0 16 0 3 1 0 0 2
144 204
144 178
1 0 2 0 0 16 0 8 0 0 11 3
52 240
52 246
143 246
2 2 3 0 0 16 0 8 7 0 0 3
52 206
52 102
121 102
1 0 2 0 0 16 0 3 0 0 15 5
144 240
144 246
143 246
143 246
220 246
1 0 5 0 0 16 0 7 0 0 13 2
144 84
144 9
2 1 5 0 0 16 0 2 5 0 0 4
105 21
105 9
220 9
220 92
3 2 7 0 0 16 0 7 1 0 0 4
144 120
144 145
144 145
144 142
1 2 2 0 0 16 0 6 5 0 0 2
220 260
220 116
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
